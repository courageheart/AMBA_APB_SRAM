///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// File Name: apb_global_pkg.sv
// Author: Farshad
// Email: farshad112@gmail.com
// Revision: 0.1
// Description: global package for holding global defines
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

package apb_global_pkg;
    // include global defines
    `include "tb_defines.sv"

endpackage